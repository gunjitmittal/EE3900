Output After Switching Initially
C1 X 0 1u ic=0
R1 X 0 1
R2 X 1 2
V2 1 0 dc 2V
.tran 100n 5u uic

.control
run
wrdata 4_7.dat v(X)
quit
.endc

.end