Amplitude Response of Butterworth Filter

V1 in 0 dc 0 ac 1
R0 in 1 1
C1 1 0 3.41m ic=0
L2 1 2 6.82m
C3 2 0 3.41m ic=0
RL 3 0 1

.control
ac dec 10 1 1000
wrdata resp_butter.txt vdb(2)
.endc

.end